library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.vga_lib.all;

-- VGA: 640x480 
-- Using the clock divider implemented in Lab 0 and your knowledge of generic component inputs, change your clock divider to accept 2 generic inputs: input frequency, and output frequency.
-- As a refresher on how the clock divider works, the clock generator should count to some value that corresponds to the number of clock pulses from the input clock there should be in the output clock
-- The output of this clock divider should be passed into the VGA entity.

-- 2. Using the provided vga_sync_gen entity, create a behavioral entity defining the behavior of the VGA synchronization signals as defined below.
-- Create two counters with equal width outputs of COUNT_RANGE as found in the provided vga_lib.vhd file.

-- h_count_r
-- Continually counts up to the horizontal period (H_MAX – See vga_lib.vhd) and then starts over at 0, using the 25 MHz pixel clock.
-- A value of zero on h_count_r corresponds to the beginning of section D in Figure 1.

-- v_count_r
-- Counts up to the vertical period (V_MAX – See vga_lib.vhd). It will increment at a particular point in the horizontal counters count (Hcount = H_VERT_INC – See vga_lib.vhd).
-- A value of zero on v_count_r corresponds to the beginning of section R in Figure 2.

-- The values of video_on, h_sync, and v_sync are determined by comparing the values of h_count_r and v_count_r with the constants provided in vga_lib.vhd

-- 3. To complete the remaining functionality of the VGA module, you will create an architecture for the provided VGA entity that instantiates the vga_sync_gen from the previous step and uses the outputs to draw a 64x64 pixel square in the center of the monitor with 12-bit hex value of #73b.

-- The VGA implementation partitions the screen into 2x2 pixel-sized blocks, each
-- of which displays a color made from a combination or red, green, and blue. There
-- will be a total of 4096 blocks arranged as a 64x64 grid, which forms a 128x128
-- image. VGA resolution is 640x480, so you must make sure the pixels not used by
-- the image are black.

-- Note that the VGA entity has a video_on output, which is not part of a normal
-- VGA interface. We are including it for verification purposes. The video_on signal
-- should connect to the video_on output of the vga_sync_gen entity. Note in the
-- top-level entity that the video_on output is left open because it is not used
-- outside of the testbench.

-- To properly determine when to draw your image, you will need to implement two
-- logical elements in your design.

-- Row bound logic: Use the v_count signal to determine the position
-- currently being drawn on the monitor. Only enable your vertical output if
-- the v_count value corresponds to the proper rows on screen.

-- Column bound logic: Use the h_count signal to determine the horizontal
-- position currently being drawn on the monitor. Only enable your horizontal
-- output if the h_count value corresponds to the proper columns on screen.

-- I recommend an enable signal that makes the color output all zero
-- if both the row and column logic don’t output one.

-- 4. Run the provided VGA testbench to test the timing of your VGA outputs and adjust your
-- timing as necessary until there are no errors remaining. This testbench will also output a
-- .txt file that can be used to simulate the VGA monitor after verifying in the testbench. It is
-- a fairly strict test for timing to make sure the outputs closely align with Figures 1, 2, & 3.

entity vga is
    port (clk              : in  std_logic;
          rst              : in  std_logic;
          en               : in  std_logic;
		  switch           : in  std_logic_vector(9 downto 0) := (others => '0');
          img_pos          : in  std_logic_vector(2 downto 0) := (others => '0');
          red, green, blue : out std_logic_vector(3 downto 0) := (others => '0');
          h_sync, v_sync   : out std_logic;
          video_on         : out std_logic);
end vga;

architecture default_arch of vga is

    signal v_count : std_logic_vector(COUNT_RANGE);
    signal h_count : std_logic_vector(COUNT_RANGE);
    -- Clocks
    signal slow_clk : std_logic := '0'; -- Slow clock
    -- Internal Temp signals
    signal temp_h_sync, temp_v_sync, temp_video_on : std_logic;
		-- x and y coordinates of ball
    signal x_pos, y_pos : integer := 200; -- 200 is the center of the screen
    signal mov_x, mov_y : integer := 1;
    -- Constants of the ball
    constant speed : integer := 2;
    constant size : integer := 64;
    constant X_MAX : integer := 638;
    constant Y_MAX : integer := 478;
    -- Constants for the paddles
    constant PADDLE_WIDTH : integer := 10;
    constant PADDLE_HEIGHT : integer := 50;
    constant PADDLE_SPEED : integer := 2;
    constant PADDLE_MAX : integer := 428;
    constant PADDLE_MIN : integer := 0;
    -- x and y coordinates for each paddle, one on the left and one on the right
    -- Paddle 1 is on the left, Paddle 2 is on the right
    signal x_pos_p1 : integer := 0;
    signal y_pos_p1 : integer := 200;
    signal x_pos_p2 : integer := 638 - PADDLE_WIDTH;
    signal y_pos_p2 : integer := 200;

    signal P1_score : integer := 0;
    signal P2_score : integer := 0;

-- BITMAPS for PONG, P1 and P2 scores, 0-9 , game over and start
-- using the 2D array to store the bitmaps
-- The dimensions of the array are 8x4
-- PONG
    type arr_type is array (0 to 7) of std_logic_vector(3 downto 0);
    type arr_type_2d is array (0 to 3, 0 to 7) of std_logic_vector(3 downto 0);
    
    signal bitmap : arr_type := ("0110", "1001", "1001", "1111", "1001", "1001", "1001", "1001");
    signal bitmap_p1 : arr_type := ("1111", "1000", "1000", "1110", "1000", "1000", "1000", "1111");
    signal bitmap_p2 : arr_type := ("1111", "0001", "0001", "0111", "0001", "0001", "0001", "1111");
    signal bitmap_0 : arr_type := ("1111", "1001", "1001", "1001", "1001", "1001", "1001", "1111");
    signal bitmap_1 : arr_type := ("0110", "0010", "0010", "0010", "0010", "0010", "0010", "1111");
    signal bitmap_2 : arr_type := ("1111", "0001", "0001", "1111", "1000", "1000", "1000", "1111");
    signal bitmap_3 : arr_type := ("1111", "0001", "0001", "0111", "0001", "0001", "0001", "1111");
    signal bitmap_4 : arr_type := ("1001", "1001", "1001", "1111", "0001", "0001", "0001", "0001");
    signal bitmap_5 : arr_type := ("1111", "1000", "1000", "1111", "0001", "0001", "0001", "1111");
    signal bitmap_6 : arr_type := ("1111", "1000", "1000", "1111", "1001", "1001", "1001", "1111");
    signal bitmap_7 : arr_type := ("1111", "0001", "0001", "0010", "0010", "0010", "0010", "0010");
    signal bitmap_8 : arr_type := ("1111", "1001", "1001", "1111", "1001", "1001", "1001", "1111");
    signal bitmap_9 : arr_type := ("1111", "1001", "1001", "1111", "0001", "0001", "0001", "1111");

    -- Position of the bitmap

    -- Position of the P1 score
    signal x_pos_p1_score : integer := 100;
    signal y_pos_p1_score : integer := 100;

    -- Position of the P2 score
    signal x_pos_p2_score : integer := 500;
    signal y_pos_p2_score : integer := 100;

begin 		
	-- Slow Clock Divider splits the 50MHz clock into 1Hz
	clk_div: entity work.clk_div
		generic map(
			clk_in_freq => 50e6,
			clk_out_freq => 20
		)
		port map(
			clk_in => clk,
			rst => rst,
			clk_out => slow_clk
		);

	-- VGA SYNC_GEN BEGINS
	sync: entity work.vga_sync_gen
		port map (clk => clk,
				    rst => rst,
				    h_count => h_count,
				    v_count => v_count,
				    h_sync => temp_h_sync,
					v_sync => temp_v_sync,
					video_on => temp_video_on);
   -- VGA_SYNC_GEN ENDS	

   -- The ball movement process
    -- The ball will move in the x and y directions
    -- The ball will bounce off top and bottom walls
    -- The ball will bounce off the paddles
    -- The ball will reset to the center of the screen it hits the left or right wall

    -- Additionally, if 'rst' is '1', the ball will reset to the center of the screen
    ball_move: process(slow_clk, rst)
        variable temp_mov_x: integer;
        variable temp_mov_y: integer;
        variable temp_x_pos: integer;
        variable temp_y_pos: integer;
    begin
        temp_mov_x := mov_x;
        temp_mov_y := mov_y;
        temp_x_pos := x_pos;
        temp_y_pos := y_pos;
        if rising_edge(slow_clk) then

            if rst = '1' then
                x_pos <= 200;
                y_pos <= 200;
                temp_mov_x := 0;
                temp_mov_y := 0;
                mov_x <= 0; -- Stopping the balls movement
                mov_y <= 0;

            else
                -- If the ball hits the left or right wall, reset the ball to the center
                if x_pos + size >= X_MAX or x_pos <= 0 then
                    -- Reset the ball to the center
                    temp_x_pos := 200;
                    temp_y_pos := 200;
                    mov_x <= 1;
                    mov_y <= 1;
                -- If the ball hits the top or bottom wall, reverse the direction of the ball
                elsif y_pos + size >= Y_MAX or y_pos <= 0 then
                    mov_y <= -1 * mov_y;
                    temp_mov_y := -1 * temp_mov_y;
                -- If the ball hits the paddle 1, reverse the direction of the ball
                elsif
                    x_pos <= x_pos_p1 + PADDLE_WIDTH and
                    y_pos + size >= y_pos_p1 and
                    y_pos <= y_pos_p1 + PADDLE_HEIGHT then
                    mov_x <= -1 * mov_x;
                    temp_mov_x := -1 * temp_mov_x;
                -- If the ball hits the paddle 2, reverse the direction of the ball
                elsif
                    x_pos + size >= x_pos_p2 and
                    y_pos + size >= y_pos_p2 and
                    y_pos <= y_pos_p2 + PADDLE_HEIGHT then
                    mov_x <= -1 * mov_x;
                    temp_mov_x := -1 * temp_mov_x;
                end if;
                x_pos <= temp_x_pos + (temp_mov_x * speed);
                y_pos <= temp_y_pos + (temp_mov_y * speed);
            end if;
        end if;
    end process ball_move;

    -- Paddle 1 movement
    -- Paddle 1 is dependent on the switches to move up and down
    -- Switches 0 and 1 are used to move the paddle up and down
    paddle1_move: process(slow_clk, rst)
        variable temp_y_pos_p1: integer;
        variable temp_x_pos_p1: integer;
    begin
        temp_y_pos_p1 := y_pos_p1;
        temp_x_pos_p1 := x_pos_p1;
        if rising_edge(slow_clk) then
            if rst = '1' then
                y_pos_p1 <= 200;
                x_pos_p1 <= 0;
            else
                if switch(0) = '1' and y_pos_p1 - PADDLE_SPEED >= PADDLE_MIN then
                    y_pos_p1 <= y_pos_p1 - PADDLE_SPEED;
                    temp_y_pos_p1 := y_pos_p1 - PADDLE_SPEED;
                elsif switch(1) = '1' and y_pos_p1 + PADDLE_SPEED <= PADDLE_MAX then
                    y_pos_p1 <= y_pos_p1 + PADDLE_SPEED;
                    temp_y_pos_p1 := y_pos_p1 + PADDLE_SPEED;
                end if;
                y_pos_p1 <= temp_y_pos_p1;
                x_pos_p1 <= temp_x_pos_p1;
            end if;
        end if;
    end process paddle1_move;

    -- Paddle 2 movement
    paddle2_move: process(slow_clk, rst)
        variable temp_y_pos_p2: integer;
        variable temp_x_pos_p2: integer;
    begin
        temp_y_pos_p2 := y_pos_p2;
        temp_x_pos_p2 := x_pos_p2;
        if rising_edge(slow_clk) then
            if rst = '1' then
                y_pos_p2 <= 200;
                x_pos_p2 <= 638 - PADDLE_WIDTH;
            else
                if switch(2) = '1' and y_pos_p2 - PADDLE_SPEED >= PADDLE_MIN then
                    y_pos_p2 <= y_pos_p2 - PADDLE_SPEED;
                    temp_y_pos_p2 := y_pos_p2 - PADDLE_SPEED;
                elsif switch(3) = '1' and y_pos_p2 + PADDLE_SPEED <= PADDLE_MAX then
                    y_pos_p2 <= y_pos_p2 + PADDLE_SPEED;
                    temp_y_pos_p2 := y_pos_p2 + PADDLE_SPEED;
                end if;
                y_pos_p2 <= temp_y_pos_p2;
                x_pos_p2 <= temp_x_pos_p2;
            end if;
        end if;
    end process paddle2_move;

	draw: process(clk, rst)
	begin
		if rising_edge(clk) then
            -- Drawing the ball
            if unsigned(h_count) >= to_unsigned(x_pos, h_count'length) and unsigned(h_count) <= to_unsigned(x_pos + size, h_count'length) and
            unsigned(v_count) >= to_unsigned(y_pos, v_count'length) and unsigned(v_count) <= to_unsigned(y_pos + size, v_count'length) and
            temp_video_on = '1' then  
                red <= "0111";
                green <= "0011";
                blue <= "1011";
            --- Paddle 1
            elsif unsigned(h_count) >= to_unsigned(x_pos_p1, h_count'length) and unsigned(h_count) <= to_unsigned(x_pos_p1 + PADDLE_WIDTH, h_count'length) and
            unsigned(v_count) >= to_unsigned(y_pos_p1, v_count'length) and unsigned(v_count) <= to_unsigned(y_pos_p1 + PADDLE_HEIGHT, v_count'length) and
            temp_video_on = '1' then
                red <= "0000";
                green <= "0000";
                blue <= "1111";
            --- Paddle 2
            elsif unsigned(h_count) >= to_unsigned(x_pos_p2, h_count'length) and unsigned(h_count) <= to_unsigned(x_pos_p2 + PADDLE_WIDTH, h_count'length) and
            unsigned(v_count) >= to_unsigned(y_pos_p2, v_count'length) and unsigned(v_count) <= to_unsigned(y_pos_p2 + PADDLE_HEIGHT, v_count'length) and
            temp_video_on = '1' then
                red <= "1111";
                green <= "0000";
                blue <= "0000";
            --- Drawing score for P1
            -- We need to draw the score and check if first we are in the display area
            -- and then check what specific pixel we are in
            -- we then check the value of the bitmap for that score at that pixel
            -- Our bitmap is 8x4 so it has 8 rows and 4 columns
            elsif unsigned(h_count) >= to_unsigned(x_pos_p1_score, h_count'length) and unsigned(h_count) <= to_unsigned(x_pos_p1_score + 4, h_count'length) and
            unsigned(v_count) >= to_unsigned(y_pos_p1_score, v_count'length) and unsigned(v_count) <= to_unsigned(y_pos_p1_score + 8, v_count'length) and
            temp_video_on = '1' then
                case P1_score is
                    when 0 =>
                        -- Draw the bitmap for 0

                        
            else
                red <= "0000";
                green <= "0000";
                blue <= "0000";
			end if;
		end if;
	end process draw;

	-- VGA MAIN ENDS
	h_sync <= temp_h_sync;
	v_sync <= temp_v_sync;
	video_on <= temp_video_on;
end default_arch;
